-- 8bit Adder
